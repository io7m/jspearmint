              