#              