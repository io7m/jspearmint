#              